TRAN RLC
*
VIN 1 0 0 PWL 0 0 10N 5
+ 25M 5 25.01M 0
L1 2 3 0.125
C1 3 0 1U
R1 1 2 200
.TRAN .2M 50M
