Alimentatore negativo
*
D1 1 3 mydiode
D2 0 2 mydiode
D3 2 3 mydiode
D4 0 1 mydiode
C 3 0 2m
RL 3 0 1k
VIN  1 2 0 AC 12 50 SIN 0 12 50
.TRAN 80m
.model mydiode D IS=10f CJ0=100F TT=100n
